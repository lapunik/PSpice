* C:\Users\Lapunik\OneDrive\Dokumenty\PSpice\ENZ\Schematic_1_cvi_Zdroj.sch

* Schematics Version 9.2
* Tue Feb 25 11:51:57 2020



** Analysis setup **
.tran 0u 100m 0 10u
.OP 


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "Schematic_1_cvi_Zdroj.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
