***E_LAPLACE_SEMESTRALKA.cir***

.LIB "nom.lib" 

.PARAM fc=2000 omega2={(2*3.1416*fc)*(2*3.1416*fc)} omega={(2*3.1416*fc)} 
.PARAM omega6={omega2*omega2*omega2}
.PARAM a1={3.588} b1={10.464} a2={0.4925} b2={1.9622} a3={0.0995} b3={1.0826}

*V1 1 0 AC 1 
V1 1 0 PULSE 0 1 1m 0 0 6m 7m
R1 1 0 1MEG 
E1 2 0 LAPLACE {V(1,0)}={(omega6/((omega2+(omega*a1*s)+(s*s*b1))*(omega2+(omega*a2*s)+(s*s*b2))*(omega2+(omega*a3*s)+(s*s*b3))))};
R2 2 0 1MEG 
.OP 
*.AC DEC 101 10 10k 
.TRAN 6u 6m 0 6u;
.PROBE V(2) 
.END
