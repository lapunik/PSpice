* C:\Users\Lapunik\OneDrive\Dokumenty\PSpice\ENZ\Schematic_1_cvi_Seriova_stabilizace_s_OZ.sch

* Schematics Version 9.2
* Tue Feb 25 12:36:42 2020


.PARAM         zatez=100 

** Analysis setup **
.DC LIN PARAM zatez 100 10m 1m 
.OP 


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "Schematic_1_cvi_Seriova_stabilizace_s_OZ.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
