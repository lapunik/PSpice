* C:\Users\Lapunik\Dropbox\PSpice\Schematics\ne5532_delic_Schematic.sch

* Schematics Version 9.2
* Thu Nov 21 12:08:37 2019



** Analysis setup **
.tran 10u 10m 0 10u
.OP 


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "C:\Users\Lapunik\Dropbox\PSpice\Knihovna_z_netu\NE5532\moje_knihovna.lib"
.lib "nom.lib"

.INC "ne5532_delic_Schematic.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
