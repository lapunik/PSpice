* C:\Users\Lapunik\Dropbox\PSpice\Schematics\Sumovy_filtr_Semestralni_prace.sch

* Schematics Version 9.2
* Wed Jan 15 08:53:23 2020


.PARAM         kondenzator35=150p 

** Analysis setup **
.ac DEC 101 100 100k
.tran 1us 2m 0 1us
.STEP  PARAM kondenzator35 LIST 
+ 100p 150p 300p
.OP 


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "C:\Users\Lapunik\Dropbox\PSpice\Knihovna_z_netu\nova\knihovna.lib"
.lib "nom.lib"

.INC "Sumovy_filtr_Semestralni_prace.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
