* C:\Users\Lapunik\Dropbox\PSpice\Schematics\Navrh_filtru_Semestralni_prace_II.sch

* Schematics Version 9.2
* Mon Dec 02 18:46:07 2019


.PARAM         odpor=1MEG 
.PARAM         fp=2 FC=1k Q=1.307

** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "C:\Users\Lapunik\Dropbox\PSpice\Knihovna_z_netu\nova\knihovna.lib"
.lib "nom.lib"

.INC "Navrh_filtru_Semestralni_prace_II.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
