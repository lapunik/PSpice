* C:\Users\Lapunik\Dropbox\PSpice\Schematics\Chyby_Druhy_Schematic.sch

* Schematics Version 9.2
* Thu Oct 10 11:43:27 2019



** Analysis setup **
.tran 10ms 10ms 0 10u
.OP 


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "Chyby_Druhy_Schematic.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
