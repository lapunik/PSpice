* C:\Users\Lapunik\Dropbox\PSpice\Schematics\statistika_schematic.sch

* Schematics Version 9.2
* Thu Nov 14 12:10:46 2019



** Analysis setup **
.ac DEC 101 10k 1MEG
.WCASE AC v([out]) YMAX
+  LIST VARY DEV LOW
.OP 


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "statistika_schematic.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
