***ne5532.cir**

.LIB "nom.lib"
.LIB "C:\Users\Lapunik\Dropbox\PSpice\Knihovna_z_netu\NE5532\moje_knihovna.lib"

*zkousime knihovnu

V1 3 0 DC 15
V2 0 4 DC 15  
V3 10 0 SIN 0 1 1k 0 0 0 
R1 10 2 1k 
R2 2 5 2k
R3 5 0 1MEG
X1 0 2 3 4 5 NE5532; volam podobvod NE5532 z knihovny

.OP
.TRAN 10u 10m 0 10u  

.PROBE V(5) V(10)

.END