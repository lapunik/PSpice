* C:\Users\Lapunik\Dropbox\PSpice\Schematics\Prvni_Schematic.sch

* Schematics Version 9.2
* Thu Oct 03 12:42:04 2019



** Analysis setup **
.tran 10u 10m 0 10u
.OP 


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "Prvni_Schematic.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
