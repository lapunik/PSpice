* C:\Users\Lapunik\Dropbox\PSpice\Schematics\VDBmarker_ schematic.sch

* Schematics Version 9.2
* Thu Oct 17 12:27:16 2019



** Analysis setup **
.ac DEC 101 10 1MEG
.tran 10u 10m 0 10u
.OP 


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "VDBmarker_ schematic.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
