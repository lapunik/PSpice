*LP_CHEBYSHEV.cir*

.LIB "nom.lib"

V1 1 0 AC 1 
R1 1 0 1MEG 
E1 2 0 CHEBYSHEV {V(1)}=LP 2k 3k 2 30 
R2 2 0 1MEG 
.OP
 
.AC DEC 101 1 100k 

.PROBE V(2) 

.END
