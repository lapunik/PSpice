* C:\Users\Lapunik\Dropbox\PSpice\Schematics\prechodak_schematic.sch

* Schematics Version 9.2
* Thu Oct 17 12:20:15 2019



** Analysis setup **
.tran 10u 10m 0 10u
.OP 


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "prechodak_schematic.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
